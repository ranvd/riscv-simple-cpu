`timescale 1ns/1ps

module rv32ima_min_sopc_tb();
    reg CLOCK_50;
    reg rst;
    
    initial begin
        CLOCK_50 = 1'b0;
        forever #10 CLOCK_50 = ~CLOCK_50;
    end
    
    inital begin
        rst = `RstEnable;
        #195 rst= `RstDisable;
        #1000 $stop;
    end
    
    rv32ima_min_sopc  rv32ima_min_sopc0(
        .clk(CLOCK_50),
        .rst(rst)
    );
endmodule