module M_extend (
    ports
);
    
endmodule